CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 311 607 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V11
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45841.8 0
0
13 Logic Switch~
5 215 607 0 1 11
0 14
0
0 0 21360 90
2 0V
14 0 28 8
3 V10
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45841.8 0
0
13 Logic Switch~
5 116 605 0 1 11
0 15
0
0 0 21360 90
2 0V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45841.8 0
0
13 Logic Switch~
5 65 416 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
45841.8 0
0
13 Logic Switch~
5 63 351 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
45841.8 0
0
13 Logic Switch~
5 63 296 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
45841.8 0
0
13 Logic Switch~
5 62 248 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
45841.8 0
0
13 Logic Switch~
5 62 195 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
45841.8 0
0
13 Logic Switch~
5 63 145 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
45841.8 0
0
13 Logic Switch~
5 62 88 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
45841.8 0
0
13 Logic Switch~
5 61 35 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
45841.8 0
0
14 Logic Display~
6 998 112 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
45841.8 0
0
5 4071~
219 862 139 0 3 22
0 4 3 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
3536 0 0
2
45841.8 0
0
8 4-In OR~
219 807 259 0 5 22
0 8 7 5 6 3
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U6B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
4597 0 0
2
45841.8 0
0
8 4-In OR~
219 632 89 0 5 22
0 12 11 10 9 4
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
3835 0 0
2
45841.8 0
0
9 Inverter~
13 397 524 0 2 22
0 13 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
3670 0 0
2
45841.8 0
0
9 Inverter~
13 281 528 0 2 22
0 14 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
5616 0 0
2
45841.8 0
0
9 Inverter~
13 170 533 0 2 22
0 15 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
9323 0 0
2
45841.8 0
0
5 4082~
219 844 508 0 5 22
0 19 15 14 13 6
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
317 0 0
2
45841.8 0
0
5 4082~
219 732 446 0 5 22
0 20 15 14 16 5
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
3108 0 0
2
45841.8 0
0
5 4082~
219 669 374 0 5 22
0 21 15 17 13 7
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
4299 0 0
2
45841.8 0
0
5 4082~
219 582 308 0 5 22
0 22 15 17 16 8
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
9672 0 0
2
45841.8 0
0
5 4082~
219 505 229 0 5 22
0 23 18 14 13 9
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
7876 0 0
2
45841.8 0
0
5 4082~
219 428 158 0 5 22
0 24 18 14 16 10
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
6369 0 0
2
45841.8 0
0
5 4082~
219 363 94 0 5 22
0 25 17 13 18 11
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
9172 0 0
2
45841.8 0
0
5 4082~
219 378 35 0 5 22
0 26 17 16 18 12
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
7100 0 0
2
45841.8 0
0
47
3 1 2 0 0 4224 0 13 12 0 0 3
895 139
998 139
998 130
5 2 3 0 0 8320 0 14 13 0 0 4
840 259
841 259
841 148
849 148
5 1 4 0 0 4224 0 15 13 0 0 4
665 89
841 89
841 130
849 130
3 5 5 0 0 8320 0 14 20 0 0 6
790 264
757 264
757 419
758 419
758 446
753 446
4 5 6 0 0 8336 0 14 19 0 0 8
790 273
794 273
794 424
880 424
880 510
866 510
866 508
865 508
2 5 7 0 0 8320 0 14 21 0 0 4
790 255
698 255
698 374
690 374
1 5 8 0 0 4224 0 14 22 0 0 4
790 246
611 246
611 308
603 308
5 4 9 0 0 8320 0 23 15 0 0 4
526 229
607 229
607 103
615 103
5 3 10 0 0 4224 0 24 15 0 0 4
449 158
602 158
602 94
615 94
5 2 11 0 0 4224 0 25 15 0 0 4
384 94
607 94
607 85
615 85
5 1 12 0 0 4224 0 26 15 0 0 4
399 35
607 35
607 76
615 76
0 4 13 0 0 4224 0 0 19 31 0 4
335 524
787 524
787 522
820 522
0 3 14 0 0 4224 0 0 19 29 0 4
234 483
792 483
792 513
820 513
0 2 15 0 0 12416 0 0 19 23 0 4
132 509
147 509
147 504
820 504
0 4 16 0 0 4096 0 0 20 34 0 2
443 460
708 460
0 3 14 0 0 0 0 0 20 29 0 2
234 451
708 451
0 2 15 0 0 0 0 0 20 23 0 2
132 442
708 442
0 4 13 0 0 0 0 0 21 31 0 4
335 389
637 389
637 388
645 388
3 0 17 0 0 4096 0 21 0 0 35 2
645 379
302 379
0 2 15 0 0 0 0 0 21 23 0 2
132 370
645 370
0 4 16 0 0 0 0 0 22 34 0 2
443 322
558 322
0 3 17 0 0 0 0 0 22 35 0 2
302 313
558 313
0 2 15 0 0 0 0 0 22 39 0 3
132 533
132 304
558 304
0 4 13 0 0 0 0 0 23 31 0 2
335 243
481 243
0 3 14 0 0 0 0 0 23 29 0 2
234 234
481 234
0 2 18 0 0 4096 0 0 23 36 0 2
201 225
481 225
0 4 16 0 0 0 0 0 24 34 0 3
390 180
390 172
404 172
0 0 16 0 0 0 0 0 0 34 34 2
372 180
381 180
3 0 14 0 0 0 0 24 0 0 38 3
404 163
234 163
234 528
0 2 18 0 0 0 0 0 24 36 0 2
201 154
404 154
3 0 13 0 0 0 0 25 0 0 37 3
339 99
335 99
335 524
0 2 17 0 0 0 0 0 25 35 0 2
302 90
339 90
0 4 18 0 0 0 0 0 25 36 0 2
201 108
339 108
2 3 16 0 0 8320 0 16 26 0 0 6
418 524
443 524
443 180
278 180
278 40
354 40
2 2 17 0 0 4224 0 17 26 0 0 5
302 528
302 58
281 58
281 31
354 31
2 4 18 0 0 8320 0 18 26 0 0 4
191 533
201 533
201 49
354 49
1 1 13 0 0 0 0 1 16 0 0 3
312 594
312 524
382 524
1 1 14 0 0 0 0 2 17 0 0 3
216 594
216 528
266 528
1 1 15 0 0 0 0 3 18 0 0 3
117 592
117 533
155 533
1 1 19 0 0 8320 0 19 4 0 0 5
820 495
820 496
86 496
86 416
77 416
1 1 20 0 0 4224 0 20 5 0 0 4
708 433
89 433
89 351
75 351
1 1 21 0 0 4224 0 21 6 0 0 4
645 361
84 361
84 296
75 296
1 1 22 0 0 4224 0 22 7 0 0 4
558 295
83 295
83 248
74 248
1 1 23 0 0 4224 0 23 8 0 0 4
481 216
83 216
83 195
74 195
1 1 24 0 0 4224 0 24 9 0 0 2
404 145
75 145
1 1 25 0 0 4224 0 25 10 0 0 4
339 81
83 81
83 88
74 88
1 1 26 0 0 4224 0 26 11 0 0 4
354 22
82 22
82 35
73 35
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
