CircuitMaker Text
5.6
Probes: 1
V5_1
Operating Point
0 429 482 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 340 30 80 10
599 88 1364 715
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.371611 0.261438
599 482 1364 715
9437202 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 195 571 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
523 0 0
2
45836.8 3
0
13 Logic Switch~
5 195 722 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6748 0 0
2
45836.8 2
0
13 Logic Switch~
5 234 632 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6901 0 0
2
45836.8 1
0
13 Logic Switch~
5 192 483 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
842 0 0
2
45836.8 0
0
7 Ground~
168 2530 710 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3277 0 0
2
45836.8 0
0
14 Logic Display~
6 2551 682 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4212 0 0
2
45836.8 0
0
14 Logic Display~
6 2541 557 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4720 0 0
2
45836.8 0
0
14 Logic Display~
6 1306 680 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5551 0 0
2
45836.8 0
0
14 Logic Display~
6 1417 722 0 1 2
10 4
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6986 0 0
2
45836.8 0
0
5 4023~
219 1578 579 0 4 22
0 6 4 4 10
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 3 6 0
1 U
8745 0 0
2
45836.8 13
0
5 4023~
219 1585 713 0 4 22
0 4 4 4 9
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 6 0
1 U
9592 0 0
2
45836.8 12
0
5 4011~
219 1734 584 0 3 22
0 10 6 4
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 7 0
1 U
8748 0 0
2
45836.8 11
0
5 4011~
219 1738 717 0 3 22
0 4 9 6
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 7 0
1 U
7168 0 0
2
45836.8 10
0
5 4011~
219 2384 703 0 3 22
0 3 7 2
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 7 0
1 U
631 0 0
2
45836.8 9
0
5 4011~
219 2380 570 0 3 22
0 8 2 3
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 7 0
1 U
9466 0 0
2
45836.8 8
0
5 4023~
219 2231 699 0 4 22
0 4 4 3 7
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 6 0
1 U
3266 0 0
2
45836.8 7
0
5 4023~
219 2224 565 0 4 22
0 2 4 4 8
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 3 5 0
1 U
7693 0 0
2
45836.8 6
0
14 Logic Display~
6 1906 699 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3723 0 0
2
45836.8 5
0
14 Logic Display~
6 1990 708 0 1 2
10 4
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3440 0 0
2
45836.8 4
0
5 4023~
219 335 574 0 4 22
0 11 18 16 15
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 5 0
1 U
6263 0 0
2
45836.8 13
0
5 4023~
219 342 708 0 4 22
0 16 17 4 14
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 5 0
1 U
4900 0 0
2
45836.8 12
0
5 4011~
219 491 579 0 3 22
0 15 11 4
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 4 0
1 U
8783 0 0
2
45836.8 11
0
5 4011~
219 495 712 0 3 22
0 4 14 11
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 4 0
1 U
3221 0 0
2
45836.8 10
0
5 4011~
219 1141 698 0 3 22
0 4 12 5
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 4 0
1 U
3215 0 0
2
45836.8 9
0
5 4011~
219 1137 565 0 3 22
0 13 5 4
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 4 0
1 U
7903 0 0
2
45836.8 8
0
5 4023~
219 988 694 0 4 22
0 4 4 4 12
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U3C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 3 3 0
1 U
7121 0 0
2
45836.8 7
0
5 4023~
219 981 560 0 4 22
0 5 4 4 13
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U3B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 3 0
1 U
4484 0 0
2
45836.8 6
0
14 Logic Display~
6 663 694 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5996 0 0
2
45836.8 5
0
14 Logic Display~
6 747 703 0 1 2
10 4
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7804 0 0
2
45836.8 4
0
57
1 0 2 0 0 4096 0 5 0 0 17 2
2530 704
2530 703
1 0 2 0 0 4096 0 6 0 0 17 2
2551 700
2551 703
1 0 3 0 0 4096 0 7 0 0 18 2
2541 575
2541 576
0 2 4 0 0 4096 0 0 17 10 0 4
1990 650
2192 650
2192 565
2200 565
1 0 5 0 0 0 0 8 0 0 39 2
1306 698
1306 698
0 0 4 0 0 0 0 0 0 31 40 2
1550 639
1417 639
0 2 4 0 0 0 0 0 11 8 0 3
1469 579
1469 713
1561 713
0 2 4 0 0 0 0 0 10 40 0 2
1417 579
1554 579
0 0 4 0 0 8320 0 0 0 31 44 3
1550 588
1550 483
846 483
0 1 4 0 0 0 0 0 19 29 0 2
1990 622
1990 694
1 0 6 0 0 4096 0 18 0 0 28 2
1906 717
1905 717
0 1 2 0 0 8320 0 0 17 17 0 5
2515 703
2515 525
2192 525
2192 556
2200 556
0 3 3 0 0 8320 0 0 16 18 0 5
2493 570
2493 723
2194 723
2194 708
2207 708
0 2 2 0 0 0 0 0 15 17 0 5
2458 703
2458 590
2348 590
2348 579
2356 579
0 1 3 0 0 0 0 0 14 18 0 5
2444 570
2444 683
2352 683
2352 694
2360 694
4 2 7 0 0 4224 0 16 14 0 0 4
2258 699
2352 699
2352 712
2360 712
3 0 2 0 0 0 0 14 0 0 0 3
2411 703
2551 703
2551 699
3 0 3 0 0 0 0 15 0 0 0 5
2407 570
2529 570
2529 576
2541 576
2541 568
4 1 8 0 0 4224 0 17 15 0 0 4
2251 565
2348 565
2348 561
2356 561
3 1 4 0 0 0 0 17 16 0 0 4
2200 574
2196 574
2196 690
2207 690
0 2 4 0 0 0 0 0 16 22 0 5
2092 622
2092 713
2199 713
2199 699
2207 699
0 0 4 0 0 16 0 0 0 9 20 6
1550 484
2091 484
2091 562
2093 562
2093 623
2196 623
0 1 6 0 0 8320 0 0 10 28 0 5
1869 717
1869 539
1546 539
1546 570
1554 570
0 3 4 0 0 0 0 0 11 29 0 5
1847 584
1847 737
1548 737
1548 722
1561 722
0 2 6 0 0 0 0 0 12 28 0 5
1812 717
1812 604
1702 604
1702 593
1710 593
0 1 4 0 0 0 0 0 13 29 0 5
1798 584
1798 697
1706 697
1706 708
1714 708
4 2 9 0 0 4224 0 11 13 0 0 4
1612 713
1706 713
1706 726
1714 726
3 0 6 0 0 0 0 13 0 0 0 3
1765 717
1905 717
1905 713
3 0 4 0 0 0 0 12 0 0 21 6
1761 584
1883 584
1883 590
1895 590
1895 622
2092 622
4 1 10 0 0 4224 0 10 12 0 0 4
1605 579
1702 579
1702 575
1710 575
3 1 4 0 0 0 0 10 11 0 0 4
1554 588
1550 588
1550 704
1561 704
0 1 4 0 0 0 0 0 29 52 0 2
747 617
747 689
1 0 11 0 0 4096 0 28 0 0 51 2
663 712
662 712
0 1 5 0 0 8320 0 0 27 39 0 5
1272 698
1272 520
949 520
949 551
957 551
0 3 4 0 0 0 0 0 26 40 0 5
1250 565
1250 718
951 718
951 703
964 703
0 2 5 0 0 0 0 0 25 39 0 5
1215 698
1215 585
1105 585
1105 574
1113 574
0 1 4 0 0 0 0 0 24 40 0 5
1201 565
1201 678
1109 678
1109 689
1117 689
4 2 12 0 0 4224 0 26 24 0 0 4
1015 694
1109 694
1109 707
1117 707
3 0 5 0 0 0 0 24 0 0 0 3
1168 698
1308 698
1308 694
3 1 4 0 0 0 0 25 9 0 0 7
1164 565
1286 565
1286 571
1298 571
1298 563
1417 563
1417 708
4 1 13 0 0 4224 0 27 25 0 0 4
1008 560
1105 560
1105 556
1113 556
3 1 4 0 0 0 0 27 26 0 0 4
957 569
953 569
953 685
964 685
0 2 4 0 0 0 0 0 26 45 0 5
849 617
849 708
956 708
956 694
964 694
1 2 4 0 0 0 0 4 27 0 0 8
204 483
848 483
848 557
853 557
853 558
949 558
949 560
957 560
0 0 4 0 0 0 0 0 0 44 42 4
848 557
849 557
849 618
953 618
0 1 11 0 0 8320 0 0 20 51 0 5
626 712
626 534
303 534
303 565
311 565
0 3 4 0 0 0 0 0 21 52 0 5
604 579
604 732
305 732
305 717
318 717
0 2 11 0 0 0 0 0 22 51 0 5
569 712
569 599
459 599
459 588
467 588
0 1 4 0 0 0 0 0 23 52 0 5
555 579
555 692
463 692
463 703
471 703
4 2 14 0 0 4224 0 21 23 0 0 4
369 708
463 708
463 721
471 721
3 0 11 0 0 0 0 23 0 0 0 3
522 712
662 712
662 708
3 0 4 0 0 0 0 22 0 0 43 6
518 579
640 579
640 585
652 585
652 617
849 617
4 1 15 0 0 4224 0 20 22 0 0 4
362 574
459 574
459 570
467 570
3 1 16 0 0 8320 0 20 21 0 0 4
311 583
307 583
307 699
318 699
1 2 17 0 0 4224 0 2 21 0 0 4
207 722
310 722
310 708
318 708
1 2 18 0 0 8320 0 1 20 0 0 5
207 571
207 572
303 572
303 574
311 574
1 0 16 0 0 0 0 3 0 0 54 2
246 632
307 632
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
