CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 370 76 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45842 0
0
13 Logic Switch~
5 213 252 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
45842 0
0
13 Logic Switch~
5 219 170 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45842 0
0
14 Logic Display~
6 572 455 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
45842 0
0
14 Logic Display~
6 574 326 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
45842 0
0
14 Logic Display~
6 573 236 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
45842 0
0
14 Logic Display~
6 578 156 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
45842 0
0
9 Inverter~
13 291 239 0 2 22
0 6 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
7361 0 0
2
45842 0
0
9 Inverter~
13 297 170 0 2 22
0 7 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
4747 0 0
2
45842 0
0
5 4073~
219 446 475 0 4 22
0 10 7 6 2
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
972 0 0
2
45842 0
0
5 4073~
219 442 350 0 4 22
0 7 10 8 3
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 1 0
1 U
3472 0 0
2
45842 0
0
5 4073~
219 439 261 0 4 22
0 10 9 6 4
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
9998 0 0
2
45842 0
0
5 4073~
219 444 174 0 4 22
0 10 9 8 5
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
3536 0 0
2
45842 0
0
18
4 1 2 0 0 4224 0 10 4 0 0 5
467 475
560 475
560 481
572 481
572 473
4 1 3 0 0 4224 0 11 5 0 0 3
463 350
574 350
574 344
4 1 4 0 0 4224 0 12 6 0 0 3
460 261
573 261
573 254
4 1 5 0 0 4224 0 13 7 0 0 5
465 174
566 174
566 182
578 182
578 174
0 3 6 0 0 4224 0 0 10 11 0 3
236 252
236 484
422 484
0 2 7 0 0 4224 0 0 10 9 0 3
262 170
262 475
422 475
0 3 8 0 0 4224 0 0 11 13 0 3
340 239
340 359
418 359
0 1 7 0 0 0 0 0 11 9 0 3
251 170
251 341
418 341
1 1 7 0 0 0 0 3 9 0 0 2
231 170
282 170
0 3 6 0 0 0 0 0 12 11 0 3
248 252
248 270
415 270
1 1 6 0 0 0 0 2 8 0 0 4
225 252
268 252
268 239
276 239
0 2 9 0 0 4096 0 0 12 14 0 3
327 170
327 261
415 261
2 3 8 0 0 0 0 8 13 0 0 4
312 239
412 239
412 183
420 183
2 2 9 0 0 4224 0 9 13 0 0 4
318 170
412 170
412 174
420 174
0 2 10 0 0 4096 0 0 11 18 0 2
370 350
418 350
0 1 10 0 0 0 0 0 12 18 0 2
370 252
415 252
0 1 10 0 0 4096 0 0 13 18 0 2
370 165
420 165
1 1 10 0 0 4224 0 1 10 0 0 3
370 88
370 466
422 466
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
