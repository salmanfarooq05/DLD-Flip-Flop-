CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 0 30 140 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 81 34 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90176e-315 0
0
13 Logic Switch~
5 200 99 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90176e-315 0
0
13 Logic Switch~
5 77 90 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90176e-315 0
0
14 Logic Display~
6 398 99 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.90176e-315 0
0
14 Logic Display~
6 575 97 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.90176e-315 0
0
14 Logic Display~
6 840 158 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.90176e-315 0
0
6 74LS76
104 644 218 0 14 29
0 6 6 4 2 2 8 9 10 11
12 5 13 14 15
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 1 0 0 0
1 U
8901 0 0
2
5.90176e-315 0
0
6 74LS76
104 452 211 0 14 29
0 6 6 3 2 2 16 17 18 19
20 4 21 22 23
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 1 0 0 0
1 U
7361 0 0
2
5.90176e-315 0
0
6 74LS76
104 286 208 0 14 29
0 6 6 7 2 2 24 25 26 27
28 3 29 30 31
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 1 0 0 0
1 U
4747 0 0
2
5.90176e-315 0
0
14 Logic Display~
6 96 380 0 1 2
10 6
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90176e-315 0
0
19
1 4 2 0 0 20608 0 1 7 0 0 8
93 34
117 34
117 39
153 39
153 34
593 34
593 209
606 209
5 0 2 0 0 0 0 9 0 0 1 3
248 208
187 208
187 34
4 0 2 0 0 0 0 9 0 0 1 3
248 199
224 199
224 34
5 0 2 0 0 0 0 8 0 0 1 3
414 211
342 211
342 34
0 4 2 0 0 0 0 0 8 1 0 3
380 34
380 202
414 202
0 5 2 0 0 0 0 0 7 1 0 3
539 34
539 218
606 218
11 1 3 0 0 4096 0 9 4 0 0 3
318 172
398 172
398 117
0 1 4 0 0 4096 0 0 5 12 0 2
575 175
575 115
11 1 5 0 0 4224 0 7 6 0 0 3
676 182
840 182
840 176
2 0 6 0 0 12416 0 7 0 0 19 4
612 191
499 191
499 309
96 309
1 0 6 0 0 0 0 7 0 0 19 4
612 182
494 182
494 288
96 288
11 3 4 0 0 4224 0 8 7 0 0 4
484 175
598 175
598 200
606 200
2 0 6 0 0 0 0 8 0 0 19 4
420 184
333 184
333 138
96 138
1 0 6 0 0 0 0 8 0 0 19 4
420 175
328 175
328 123
96 123
11 3 3 0 0 4224 0 9 8 0 0 4
318 172
406 172
406 193
414 193
1 3 7 0 0 8320 0 2 9 0 0 4
212 99
240 99
240 190
248 190
2 0 6 0 0 0 0 9 0 0 19 2
254 181
96 181
1 0 6 0 0 0 0 9 0 0 19 2
254 172
96 172
1 1 6 0 0 0 0 3 10 0 0 3
89 90
96 90
96 366
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
