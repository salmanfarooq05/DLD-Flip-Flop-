CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 607 49 0 1 11
0 5
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45841.9 0
0
13 Logic Switch~
5 528 50 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45841.9 0
0
13 Logic Switch~
5 457 52 0 1 11
0 6
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45841.9 0
0
13 Logic Switch~
5 376 55 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
45841.9 0
0
13 Logic Switch~
5 300 57 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8157 0 0
2
45841.9 0
0
13 Logic Switch~
5 231 61 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5572 0 0
2
45841.9 0
0
13 Logic Switch~
5 177 62 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8901 0 0
2
45841.9 0
0
13 Logic Switch~
5 116 65 0 1 11
0 12
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
45841.9 0
0
14 Logic Display~
6 870 317 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
45841.9 0
0
14 Logic Display~
6 870 210 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
45841.9 0
0
14 Logic Display~
6 871 85 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
45841.9 0
0
8 4-In OR~
219 737 333 0 5 22
0 8 7 6 5 2
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
9998 0 0
2
45841.9 0
0
8 4-In OR~
219 737 223 0 5 22
0 10 7 9 5 3
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U1B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
3536 0 0
2
45841.9 0
0
8 4-In OR~
219 737 111 0 5 22
0 11 6 5 9 4
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
4597 0 0
2
45841.9 0
0
14 Logic Display~
6 606 527 0 1 2
10 5
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L8
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
45841.9 0
0
14 Logic Display~
6 527 528 0 1 2
10 9
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L7
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
45841.9 0
0
14 Logic Display~
6 456 531 0 1 2
10 6
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
45841.9 0
0
14 Logic Display~
6 376 531 0 1 2
10 11
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9323 0 0
2
45841.9 0
0
14 Logic Display~
6 301 524 0 1 2
10 7
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
317 0 0
2
45841.9 0
0
14 Logic Display~
6 231 528 0 1 2
10 10
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
45841.9 0
0
14 Logic Display~
6 177 528 0 1 2
10 8
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
45841.9 0
0
14 Logic Display~
6 116 525 0 1 2
10 12
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
45841.9 0
0
23
1 5 2 0 0 8320 0 9 12 0 0 5
870 335
870 339
778 339
778 333
770 333
1 5 3 0 0 8320 0 10 13 0 0 5
870 228
870 232
778 232
778 223
770 223
5 1 4 0 0 4224 0 14 11 0 0 3
770 111
871 111
871 103
4 0 5 0 0 4096 0 12 0 0 16 2
720 347
607 347
3 0 6 0 0 4096 0 12 0 0 18 2
720 338
457 338
2 0 7 0 0 4096 0 12 0 0 20 2
720 329
300 329
1 0 8 0 0 4224 0 12 0 0 22 2
720 320
177 320
4 0 5 0 0 0 0 13 0 0 16 4
720 237
612 237
612 238
607 238
3 0 9 0 0 4096 0 13 0 0 17 2
720 228
528 228
2 0 7 0 0 0 0 13 0 0 20 4
720 219
305 219
305 220
300 220
1 0 10 0 0 4224 0 13 0 0 21 2
720 210
231 210
3 0 5 0 0 0 0 14 0 0 16 2
720 116
607 116
0 4 9 0 0 0 0 0 14 17 0 2
528 125
720 125
0 2 6 0 0 0 0 0 14 18 0 4
457 108
712 108
712 107
720 107
0 1 11 0 0 4096 0 0 14 19 0 2
376 98
720 98
1 1 5 0 0 4224 0 1 15 0 0 4
607 61
607 507
606 507
606 513
1 1 9 0 0 4224 0 2 16 0 0 3
528 62
528 514
527 514
1 1 6 0 0 4224 0 3 17 0 0 4
457 64
457 511
456 511
456 517
1 1 11 0 0 4224 0 4 18 0 0 2
376 67
376 517
1 1 7 0 0 4224 0 5 19 0 0 4
300 69
300 506
301 506
301 510
1 1 10 0 0 0 0 6 20 0 0 2
231 73
231 514
1 1 8 0 0 0 0 7 21 0 0 2
177 74
177 514
1 1 12 0 0 4224 0 8 22 0 0 2
116 77
116 511
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
