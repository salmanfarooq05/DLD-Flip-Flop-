CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 404 192 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45841.2 11
0
13 Logic Switch~
5 344 190 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45841.2 10
0
13 Logic Switch~
5 286 189 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45841.2 9
0
13 Logic Switch~
5 121 193 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
45841.2 8
0
13 Logic Switch~
5 179 194 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
45841.2 7
0
13 Logic Switch~
5 239 196 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
45841.2 6
0
13 Logic Switch~
5 472 103 0 1 11
0 20
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
45841.2 2
0
14 Logic Display~
6 1200 132 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
45841.2 0
0
14 Logic Display~
6 1170 492 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
45841.2 0
0
14 Logic Display~
6 820 174 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
45841.2 0
0
14 Logic Display~
6 710 176 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
45841.2 0
0
8 2-In OR~
219 1178 279 0 3 22
0 7 6 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9998 0 0
2
45841.2 0
0
9 2-In AND~
219 1098 244 0 3 22
0 9 8 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3536 0 0
2
45841.2 0
0
9 2-In AND~
219 1108 327 0 3 22
0 11 10 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
4597 0 0
2
45841.2 0
0
9 2-In XOR~
219 1039 435 0 3 22
0 11 10 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3835 0 0
2
45841.2 0
0
9 2-In XOR~
219 964 375 0 3 22
0 9 8 11
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3670 0 0
2
45841.2 0
0
8 2-In OR~
219 822 494 0 3 22
0 13 12 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5616 0 0
2
45841.2 0
0
9 2-In AND~
219 731 540 0 3 22
0 15 14 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9323 0 0
2
45841.2 0
0
9 2-In AND~
219 733 453 0 3 22
0 17 16 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
317 0 0
2
45841.2 0
0
9 2-In XOR~
219 751 298 0 3 22
0 17 16 4
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3108 0 0
2
45841.2 0
0
9 2-In XOR~
219 659 387 0 3 22
0 15 14 17
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4299 0 0
2
45841.2 0
0
9 2-In AND~
219 529 344 0 3 22
0 19 18 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9672 0 0
2
45841.2 0
0
14 Logic Display~
6 406 493 0 1 2
10 19
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
45841.2 14
0
14 Logic Display~
6 346 491 0 1 2
10 15
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6369 0 0
2
45841.2 13
0
14 Logic Display~
6 288 491 0 1 2
10 9
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9172 0 0
2
45841.2 12
0
14 Logic Display~
6 123 495 0 1 2
10 8
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7100 0 0
2
45841.2 5
0
14 Logic Display~
6 181 495 0 1 2
10 14
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3820 0 0
2
45841.2 4
0
14 Logic Display~
6 241 497 0 1 2
10 18
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7678 0 0
2
45841.2 3
0
9 2-In XOR~
219 534 232 0 3 22
0 19 18 21
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
961 0 0
2
45841.2 1
0
9 2-In XOR~
219 615 276 0 3 22
0 21 20 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3178 0 0
2
45841.2 0
0
36
1 3 2 0 0 4224 0 8 12 0 0 5
1200 150
1200 260
1219 260
1219 279
1211 279
3 1 3 0 0 4224 0 15 9 0 0 5
1072 435
1157 435
1157 518
1170 518
1170 510
1 3 4 0 0 4224 0 10 20 0 0 3
820 192
820 298
784 298
1 3 5 0 0 4224 0 11 30 0 0 3
710 194
710 276
648 276
3 2 6 0 0 8320 0 14 12 0 0 4
1129 327
1157 327
1157 288
1165 288
3 1 7 0 0 4224 0 13 12 0 0 4
1119 244
1157 244
1157 270
1165 270
0 2 8 0 0 8192 0 0 13 13 0 3
847 407
847 253
1074 253
0 1 9 0 0 8192 0 0 13 14 0 3
843 366
843 235
1074 235
0 2 10 0 0 8320 0 0 14 11 0 3
915 494
915 336
1084 336
0 1 11 0 0 8320 0 0 14 12 0 3
1015 375
1015 318
1084 318
3 2 10 0 0 0 0 17 15 0 0 4
855 494
1015 494
1015 444
1023 444
3 1 11 0 0 0 0 16 15 0 0 4
997 375
1015 375
1015 426
1023 426
0 2 8 0 0 4224 0 0 16 33 0 4
121 407
940 407
940 384
948 384
0 1 9 0 0 4224 0 0 16 36 0 2
286 366
948 366
3 2 12 0 0 4224 0 18 17 0 0 4
752 540
801 540
801 503
809 503
3 1 13 0 0 4224 0 19 17 0 0 4
754 453
801 453
801 485
809 485
0 2 14 0 0 4224 0 0 18 32 0 4
179 427
694 427
694 549
707 549
1 0 15 0 0 4224 0 18 0 0 35 4
707 531
359 531
359 414
344 414
0 2 16 0 0 8192 0 0 19 21 0 3
578 344
578 462
709 462
0 1 17 0 0 4096 0 0 19 22 0 3
701 387
701 444
709 444
3 2 16 0 0 4224 0 22 20 0 0 4
550 344
715 344
715 307
735 307
3 1 17 0 0 8320 0 21 20 0 0 4
692 387
720 387
720 289
735 289
0 2 14 0 0 0 0 0 21 32 0 2
179 396
643 396
0 1 15 0 0 0 0 0 21 35 0 2
344 378
643 378
0 2 18 0 0 4096 0 0 22 31 0 2
239 353
505 353
0 1 19 0 0 4096 0 0 22 34 0 2
404 335
505 335
1 2 20 0 0 4224 0 7 30 0 0 3
472 115
472 285
599 285
3 1 21 0 0 8320 0 29 30 0 0 4
567 232
591 232
591 267
599 267
0 2 18 0 0 4224 0 0 29 31 0 2
239 241
518 241
0 1 19 0 0 4096 0 0 29 34 0 2
404 223
518 223
1 1 18 0 0 0 0 6 28 0 0 4
239 208
239 478
241 478
241 483
1 1 14 0 0 0 0 5 27 0 0 4
179 206
179 476
181 476
181 481
1 1 8 0 0 0 0 4 26 0 0 4
121 205
121 475
123 475
123 481
1 1 19 0 0 4224 0 1 23 0 0 4
404 204
404 474
406 474
406 479
1 1 15 0 0 0 0 2 24 0 0 4
344 202
344 472
346 472
346 477
1 1 9 0 0 0 0 3 25 0 0 4
286 201
286 471
288 471
288 477
13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1206 250 1241 272
1215 257 1231 273
2 C2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1065 401 1102 423
1075 408 1091 424
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
849 466 884 488
858 474 874 490
2 C1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
779 266 814 288
788 274 804 290
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
546 315 581 337
555 323 571 339
2 C0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
640 244 675 266
649 251 665 267
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
451 37 494 59
460 44 484 60
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
394 122 429 143
403 129 419 144
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
332 123 365 144
340 129 356 144
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
274 126 309 147
283 133 299 148
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
229 126 264 147
238 133 254 148
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
167 127 200 148
175 134 191 149
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
109 130 144 151
118 137 134 152
2 B2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
