CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 70 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 478 122 0 1 11
0 11
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6369 0 0
2
5.90173e-315 0
0
13 Logic Switch~
5 370 125 0 1 11
0 12
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
5.90173e-315 0
0
13 Logic Switch~
5 265 128 0 1 11
0 13
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7100 0 0
2
5.90173e-315 0
0
13 Logic Switch~
5 170 289 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
5.90173e-315 0
0
14 Logic Display~
6 767 891 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.90173e-315 0
0
14 Logic Display~
6 772 814 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90173e-315 0
0
14 Logic Display~
6 776 722 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.90173e-315 0
0
14 Logic Display~
6 777 637 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.90173e-315 0
0
14 Logic Display~
6 779 548 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.90173e-315 0
0
14 Logic Display~
6 782 461 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.90173e-315 0
0
14 Logic Display~
6 782 377 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.90173e-315 0
0
14 Logic Display~
6 781 296 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
5.90173e-315 0
0
5 4082~
219 588 900 0 5 22
0 13 12 11 10 2
0
0 0 608 0
4 4082
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
9442 0 0
2
5.90173e-315 0
0
5 4082~
219 588 823 0 5 22
0 13 12 14 10 3
0
0 0 608 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
9424 0 0
2
5.90173e-315 0
0
5 4082~
219 590 732 0 5 22
0 13 15 11 10 4
0
0 0 608 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
9968 0 0
2
5.90173e-315 0
0
5 4082~
219 592 646 0 5 22
0 13 15 14 10 5
0
0 0 608 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
9281 0 0
2
5.90173e-315 0
0
5 4082~
219 592 557 0 5 22
0 16 12 11 10 6
0
0 0 608 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
8464 0 0
2
5.90173e-315 0
0
5 4082~
219 595 470 0 5 22
0 16 12 14 10 7
0
0 0 608 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
7168 0 0
2
5.90173e-315 0
0
5 4082~
219 595 386 0 5 22
0 16 15 11 10 8
0
0 0 608 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
3171 0 0
2
5.90173e-315 0
0
5 4082~
219 594 305 0 5 22
0 14 15 16 10 9
0
0 0 608 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
4139 0 0
2
5.90173e-315 0
0
9 Inverter~
13 475 209 0 2 22
0 11 14
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
6435 0 0
2
5.90173e-315 0
0
9 Inverter~
13 367 209 0 2 22
0 12 15
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
5283 0 0
2
5.90173e-315 0
0
9 Inverter~
13 262 214 0 2 22
0 13 16
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6874 0 0
2
5.90173e-315 0
0
44
5 0 2 0 0 0 0 13 0 0 2 2
609 900
609 900
5 1 2 0 0 4224 0 0 5 0 0 5
601 900
755 900
755 917
767 917
767 909
1 5 3 0 0 16512 0 6 14 0 0 5
772 832
772 840
760 840
760 823
609 823
5 1 4 0 0 8320 0 15 7 0 0 6
611 732
611 731
764 731
764 748
776 748
776 740
5 1 5 0 0 4224 0 16 8 0 0 5
613 646
765 646
765 663
777 663
777 655
5 1 6 0 0 4224 0 17 9 0 0 5
613 557
767 557
767 574
779 574
779 566
5 1 7 0 0 4224 0 18 10 0 0 5
616 470
770 470
770 487
782 487
782 479
5 1 8 0 0 4224 0 19 11 0 0 5
616 386
770 386
770 403
782 403
782 395
5 1 9 0 0 4224 0 20 12 0 0 5
615 305
769 305
769 322
781 322
781 314
4 0 10 0 0 4096 0 14 0 0 17 2
564 837
199 837
4 0 10 0 0 4096 0 15 0 0 17 2
566 746
199 746
4 0 10 0 0 4096 0 16 0 0 17 2
568 660
199 660
4 0 10 0 0 0 0 17 0 0 17 2
568 571
199 571
4 0 10 0 0 4096 0 18 0 0 17 2
571 484
199 484
0 4 10 0 0 0 0 0 19 17 0 2
199 400
571 400
0 4 10 0 0 0 0 0 20 17 0 2
199 319
570 319
1 4 10 0 0 8320 0 4 13 0 0 4
182 289
199 289
199 914
564 914
0 3 11 0 0 4096 0 0 13 24 0 3
435 736
435 905
564 905
0 2 12 0 0 8192 0 0 13 22 0 3
342 819
342 896
564 896
0 1 13 0 0 12288 0 0 13 23 0 4
300 809
303 809
303 887
564 887
0 3 14 0 0 8192 0 0 14 27 0 4
459 651
460 651
460 828
564 828
0 2 12 0 0 4096 0 0 14 31 0 3
339 553
339 819
564 819
0 1 13 0 0 8192 0 0 14 26 0 3
300 719
300 810
564 810
0 3 11 0 0 4096 0 0 15 30 0 3
435 561
435 737
566 737
0 2 15 0 0 12288 0 0 15 28 0 4
372 642
373 642
373 728
566 728
0 1 13 0 0 12288 0 0 15 29 0 4
236 633
295 633
295 719
566 719
0 3 14 0 0 0 0 0 16 33 0 4
460 475
459 475
459 651
568 651
0 2 15 0 0 8320 0 0 16 37 0 4
371 381
372 381
372 642
568 642
0 1 13 0 0 8320 0 0 16 44 0 4
265 182
236 182
236 633
568 633
0 3 11 0 0 0 0 0 17 36 0 3
435 391
435 562
568 562
0 2 12 0 0 0 0 0 17 34 0 3
336 466
336 553
568 553
0 1 16 0 0 8192 0 0 17 35 0 3
267 457
267 544
568 544
0 3 14 0 0 8320 0 0 18 41 0 4
478 292
460 292
460 475
571 475
0 2 12 0 0 8320 0 0 18 43 0 4
370 173
336 173
336 466
571 466
0 1 16 0 0 12416 0 0 18 38 0 4
268 370
264 370
264 457
571 457
0 3 11 0 0 8320 0 0 19 42 0 4
478 173
435 173
435 391
571 391
0 2 15 0 0 0 0 0 19 40 0 4
370 298
371 298
371 382
571 382
0 1 16 0 0 0 0 0 19 39 0 3
268 310
268 373
571 373
2 3 16 0 0 0 0 23 20 0 0 3
265 232
265 310
570 310
2 2 15 0 0 0 0 22 20 0 0 3
370 227
370 301
570 301
2 1 14 0 0 0 0 21 20 0 0 3
478 227
478 292
570 292
1 1 11 0 0 0 0 1 21 0 0 2
478 134
478 191
1 1 12 0 0 0 0 2 22 0 0 2
370 137
370 191
1 1 13 0 0 0 0 3 23 0 0 2
265 140
265 196
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
