CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 0 30 200 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 114 275 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45841.5 0
0
13 Logic Switch~
5 138 28 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45841.5 0
0
13 Logic Switch~
5 134 100 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
45841.5 0
0
9 Inverter~
13 173 28 0 2 22
0 4 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3421 0 0
2
45841.5 0
0
14 Logic Display~
6 638 63 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
45841.5 0
0
14 Logic Display~
6 425 57 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
45841.5 0
0
14 Logic Display~
6 320 62 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
45841.5 0
0
9 2-In AND~
219 476 117 0 3 22
0 7 6 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7361 0 0
2
45841.5 0
0
6 74LS76
104 559 201 0 14 29
0 8 8 3 2 2 10 11 12 13
14 5 15 16 17
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
4747 0 0
2
45841.5 0
0
6 74LS76
104 414 200 0 14 29
0 7 7 3 2 2 18 19 20 21
22 6 23 24 25
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
972 0 0
2
45841.5 0
0
6 74LS76
104 267 195 0 14 29
0 9 9 3 2 2 26 27 28 29
30 7 31 32 33
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
3472 0 0
2
45841.5 0
0
21
0 0 2 0 0 4096 0 0 0 6 3 2
217 195
217 275
0 0 2 0 0 0 0 0 0 5 3 2
365 200
365 275
1 0 2 0 0 4224 0 1 0 0 4 3
126 275
510 275
510 201
4 5 2 0 0 16 0 9 9 0 0 4
521 192
496 192
496 201
521 201
4 5 2 0 0 0 0 10 10 0 0 4
376 191
358 191
358 200
376 200
4 5 2 0 0 0 0 11 11 0 0 4
229 186
210 186
210 195
229 195
2 3 3 0 0 4224 0 4 9 0 0 4
194 28
513 28
513 183
521 183
0 3 3 0 0 0 0 0 11 7 0 3
210 28
210 177
229 177
0 3 3 0 0 0 0 0 10 7 0 3
369 28
369 182
376 182
1 1 4 0 0 4224 0 2 4 0 0 2
150 28
158 28
1 11 5 0 0 4224 0 5 9 0 0 3
638 81
638 165
591 165
1 0 6 0 0 4224 0 6 0 0 16 4
425 75
425 145
449 145
449 164
0 1 7 0 0 4096 0 0 7 18 0 2
320 159
320 80
3 0 8 0 0 8320 0 8 0 0 17 4
497 117
499 117
499 171
502 171
0 1 7 0 0 8320 0 0 8 18 0 3
324 159
324 108
452 108
11 2 6 0 0 0 0 10 8 0 0 4
446 164
453 164
453 126
452 126
1 2 8 0 0 0 0 9 9 0 0 4
527 165
502 165
502 174
527 174
11 0 7 0 0 0 0 11 0 0 19 4
299 159
358 159
358 169
363 169
1 2 7 0 0 0 0 10 10 0 0 4
382 164
363 164
363 173
382 173
1 0 9 0 0 8320 0 3 0 0 21 4
146 100
188 100
188 163
193 163
1 2 9 0 0 0 0 11 11 0 0 4
235 159
193 159
193 168
235 168
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
