CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
650 150 30 150 10
223 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
391 176 504 273
9437202 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 862 241 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3178 0 0
2
45841.5 2
0
13 Logic Switch~
5 862 421 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3409 0 0
2
45841.5 1
0
13 Logic Switch~
5 857 319 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3951 0 0
2
45841.5 0
0
13 Logic Switch~
5 32 327 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
45841.5 0
0
13 Logic Switch~
5 37 429 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3780 0 0
2
45841.5 0
0
13 Logic Switch~
5 37 249 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9265 0 0
2
45841.5 0
0
6 74LS76
104 1019 324 0 14 29
0 16 16 14 15 15 49 50 51 52
53 13 54 55 56
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U6
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
9442 0 0
2
45841.5 8
0
6 74LS76
104 1203 324 0 14 29
0 16 16 13 15 15 57 58 59 60
61 12 62 63 64
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
9424 0 0
2
45841.5 7
0
6 74LS76
104 1384 324 0 14 29
0 16 16 12 15 15 65 66 67 68
69 11 70 71 72
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
9968 0 0
2
45841.5 6
0
14 Logic Display~
6 1108 355 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9281 0 0
2
45841.5 5
0
14 Logic Display~
6 1300 367 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8464 0 0
2
45841.5 4
0
14 Logic Display~
6 1494 363 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
45841.5 3
0
14 Logic Display~
6 669 371 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3171 0 0
2
45841.5 0
0
14 Logic Display~
6 475 375 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4139 0 0
2
45841.5 0
0
14 Logic Display~
6 283 363 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6435 0 0
2
45841.5 0
0
6 74LS76
104 559 332 0 14 29
0 24 24 20 23 23 73 74 75 76
77 78 17 79 80
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
5283 0 0
2
45841.5 0
0
6 74LS76
104 378 332 0 14 29
0 24 24 21 23 23 81 82 83 84
85 20 18 86 87
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
6874 0 0
2
45841.5 0
0
6 74LS76
104 194 332 0 14 29
0 24 24 22 23 23 88 89 90 91
92 21 19 93 94
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
5305 0 0
2
45841.5 0
0
36
11 1 11 0 0 8320 0 9 12 0 0 5
1416 288
1481 288
1481 389
1494 389
1494 381
0 1 12 0 0 4224 0 0 11 4 0 4
1262 288
1262 393
1300 393
1300 385
0 1 13 0 0 4224 0 0 10 5 0 4
1075 277
1075 381
1108 381
1108 373
11 3 12 0 0 0 0 8 9 0 0 4
1235 288
1278 288
1278 306
1346 306
11 3 13 0 0 0 0 7 8 0 0 5
1051 288
1051 277
1101 277
1101 306
1165 306
1 3 14 0 0 8320 0 3 7 0 0 3
869 319
869 306
981 306
0 0 15 0 0 4096 0 0 0 12 9 2
962 324
962 421
0 0 15 0 0 0 0 0 0 11 9 2
1152 324
1152 421
1 0 15 0 0 4224 0 2 0 0 10 3
874 421
1335 421
1335 324
4 5 15 0 0 0 0 9 9 0 0 4
1346 315
1315 315
1315 324
1346 324
4 5 15 0 0 0 0 8 8 0 0 4
1165 315
1139 315
1139 324
1165 324
4 5 15 0 0 0 0 7 7 0 0 4
981 315
947 315
947 324
981 324
0 0 16 0 0 4096 0 0 0 15 16 2
962 241
962 288
0 0 16 0 0 0 0 0 0 15 17 2
1155 241
1155 288
1 0 16 0 0 4224 0 1 0 0 18 3
874 241
1331 241
1331 288
1 2 16 0 0 0 0 7 7 0 0 4
987 288
947 288
947 297
987 297
1 2 16 0 0 0 0 8 8 0 0 4
1171 288
1140 288
1140 297
1171 297
1 2 16 0 0 0 0 9 9 0 0 4
1352 288
1312 288
1312 297
1352 297
12 1 17 0 0 8320 0 16 13 0 0 5
597 305
656 305
656 397
669 397
669 389
12 1 18 0 0 8320 0 17 14 0 0 5
416 305
442 305
442 401
475 401
475 393
12 1 19 0 0 8320 0 18 15 0 0 5
232 305
270 305
270 389
283 389
283 381
11 3 20 0 0 12416 0 17 16 0 0 4
410 296
453 296
453 314
521 314
11 3 21 0 0 16512 0 18 17 0 0 5
226 296
226 285
276 285
276 314
340 314
1 3 22 0 0 8320 0 4 18 0 0 3
44 327
44 314
156 314
0 0 23 0 0 4096 0 0 0 30 27 2
137 332
137 429
0 0 23 0 0 0 0 0 0 29 27 2
327 332
327 429
1 0 23 0 0 4224 0 5 0 0 28 3
49 429
510 429
510 332
4 5 23 0 0 0 0 16 16 0 0 4
521 323
490 323
490 332
521 332
4 5 23 0 0 0 0 17 17 0 0 4
340 323
314 323
314 332
340 332
4 5 23 0 0 0 0 18 18 0 0 4
156 323
122 323
122 332
156 332
0 0 24 0 0 4096 0 0 0 33 34 2
137 249
137 296
0 0 24 0 0 0 0 0 0 33 35 2
330 249
330 296
1 0 24 0 0 4224 0 6 0 0 36 3
49 249
506 249
506 296
1 2 24 0 0 0 0 18 18 0 0 4
162 296
122 296
122 305
162 305
1 2 24 0 0 0 0 17 17 0 0 4
346 296
315 296
315 305
346 305
1 2 24 0 0 0 0 16 16 0 0 4
527 296
487 296
487 305
527 305
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 28
1086 507 1325 531
1093 513 1317 529
28 3 bit Asynchronus up counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
877 211 940 235
884 217 932 233
6 Inputs
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
869 281 908 305
876 286 900 302
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
864 420 951 444
871 426 943 442
9 Set Reset
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
39 428 126 452
46 434 118 450
9 Set Reset
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
44 289 83 313
51 294 75 310
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
52 219 115 243
59 225 107 241
6 Inputs
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 30
261 515 516 539
268 521 508 537
30 3 bit Asynchronus down counter
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
